module change_machine(
    input logic [3:0] cost, paid,
    input logic [1:0] quarters, dimes,nickles
    output logic [2:0] first_coin, second_coin,
    output logic exact_amount, cough_up_more, 
    output logic [3:0] remaining 
);

endmodule