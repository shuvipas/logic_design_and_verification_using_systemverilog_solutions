module p3_4 (
    input logic x,clk, rst,
    output logic y,z 
);

endmodule